----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:16:23 04/07/2021 
-- Design Name: 
-- Module Name:    adder_plus4_incrementor - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity adder_plus4_incrementor is
		Port ( input : in  STD_LOGIC_vector(31 downto 0);
             output : out  STD_LOGIC_vector(31 downto 0)
			  );
end adder_plus4_incrementor;

architecture Behavioral of adder_plus4_incrementor is
	signal inter_out : signed(31 downto 0);
	
begin 
	
	inter_out <= signed(input) + 4;
	output <= std_logic_vector(inter_out);
	
end Behavioral;


